module halfadder(s,c,a,b);
    input a,b;
    output s,c;
endmodule